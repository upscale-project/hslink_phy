/****************************************************************

Copyright (c) #YEAR# #LICENSOR#. All rights reserved.

The information and source code contained herein is the 
property of #LICENSOR#, and may not be disclosed or
reproduced in whole or in part without explicit written 
authorization from #LICENSOR#.

* Filename   : adc_clkgen.sv
* Author     : Byongchan Lim (bclim@stanford.edu)
* Description: Generate multi-phase clocks for TI-ADC
  - The input clock source is a high-speed, PI-controlled
    clock, the clock rate depends on 'Nti':
    - Nti == 1: running at full-rate ( 5.0 GHz for 5 Gbps link)
    - Nti != 1: running at half-rate ( 2.5 GHz for 5 Gbps link)
  - When Nti != 1, Nti must be multiples of 4.

* Note       :
  - If 'Nti'==1, it is non-TI-ADC configuration.
  - TI hierarchy is assumed to be Nbr x Nleaf where Nbr is
    the number of branches and Nleaf is the number of leaves 
    per branch.  This means that Nbr x Nleaf is the total number 
    of time-interleaving slices.
  - For now, Nbr is fixed to 4.

          |---
    |-----|---
    |     | .
    |     |---
    |
  --|
    |     |---
    |-----|---
    |     | .
    |     |---
    |
           ...

    Nbr     Nleaf

* Todo       :
  -

* Revision   :
  - 00/00/00: Initial commit

****************************************************************/


module adc_clkgen #(
// parameters here
  parameter integer Nti = 1 // total number of slices
) (
// I/Os here
  input cki,  // full(half)-rate clock input
  output [3:0] cko_ti_iq, // I/Q clocks for branch switch controls
                          // valid only when (Nti != 1)
  output [Nti-1:0] cko_ti_leaf // sampling clock for leaf S/H
                               // outputs in sequence from 0 to Nti-1
);

`get_timeunit

///////////////////
// CODE STARTS HERE
///////////////////

//----- SIGNAL DECLARATION -----
localparam integer Nleaf = (Nti >> 2); // number of leaves per branch
localparam [Nleaf-1:0] ck_leaf_init = {{(Nleaf-1){1'b0}}, 1'b1};
localparam logic cfg_ti = (Nti != 1);

genvar i;
logic [Nleaf-1:0] _cko_ti_leaf[3:0];

// Nti must be multiples of 4
initial 
  if (cfg_ti) assert (Nti == 4*Nleaf) else $warning("[%m:] Nti (%d) != 4*Nleaf (%d) ", Nti, 4*Nleaf);

//----- FUNCTIONAL DESCRIPTION -----
`protect
//pragma protect 
//pragma protect begin

`generate_random_seed(1,0)
real tskew[Nti];
initial begin
  for (int i=0;i<Nti;i++) tskew[i] = $dist_uniform(seed, 1, 20)*1e-12;
end

clk_iq_div iCLKGEN_IQ ( .cki(cki), .rstn(cfg_ti), .cko(cko_ti_iq) ); 

// multi-phase clocks generated by I-clock
clkgen_mph #( .Np(Nleaf), .init(ck_leaf_init) ) iCLKGEN_MPH_ ( .cki(cko_ti_iq[0]), .cko(_cko_ti_leaf[0]) );
generate

  for (i=1;i<4;i++) begin : iCLKGEN_MPH // generate rest of ti-adc clocks
    if (Nleaf == 1)
      assign _cko_ti_leaf[i] = cko_ti_iq[i];
    else
      always @(posedge cko_ti_iq[i]) _cko_ti_leaf[i] <= _cko_ti_leaf[i-1];
  end

  for (i=0;i<Nti;i++) begin : iCLKASGN  // rearrange the index of multi-phase clocks
    //assign `delay(tskew[i]) cko_ti_leaf[i] = cfg_ti ? _cko_ti_leaf[i%4][i/4] : cki;
    assign cko_ti_leaf[i] = cfg_ti ? _cko_ti_leaf[i%4][i/4] : cki;
  end

endgenerate

//pragma protect end
`endprotect

endmodule

